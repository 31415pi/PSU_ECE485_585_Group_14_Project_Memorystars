`ifdef SHOW_ALL
`define SHOW_INFILE
`define SHOW_FILENAME
`define SHOW_READ
`define SHOW_OPEN
`endif
module tb_top;
  parser tf_parser();
  
endmodule
