module tb_top;
  `timescale 1fs/1fs
  parser parsing();

endmodule
