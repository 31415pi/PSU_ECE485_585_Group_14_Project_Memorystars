module tb_top;
  `timescale 1fs/1fs
//  input logic [2:0]clk_ensig,
  parser parsing
  ();
  //  initial begin
  //  $display("tb instantiation");
//  mc mcc(
  //  .clk_en(),
   // .request(),
   // .clock(),
   // .parser_dr(),
   // .new_instruction()
 // );// tf_parser();
  // end

endmodule
